----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 	Fernando Candelario Herrero
-- Create Date:    12:19:20 05/22/2018 
-- Design Name: 
-- Module Name:    vgaTecladoInterface - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity vgaTecladoInterface is
port(
    rst_n    	: in    std_logic;
    clk        : in    std_logic;
	 teclaPulsada : in  std_logic_vector(24 downto 0);
	 hSync   	: out std_logic;
    vSync   	: out std_logic;
    RGB     	: out std_logic_vector(8 downto 0)
 );
end vgaTecladoInterface;

library ieee, unisim;
use ieee.numeric_std.all;
use unisim.vcomponents.all;
use work.common.all;

architecture Behavioral of vgaTecladoInterface is
	
	signal Pentagramas, Teclas, colorVerde, colorAzul, Notas: std_logic;
	
	signal nota : std_logic_vector(14 downto 0);
	signal teclaPulsadaPintar, notaPintar : std_logic_vector(24 downto 0);
	signal lineAux, pixelAux : std_logic_vector(9 downto 0);
	
	signal dir : std_logic_vector(8 downto 0);

	signal pixel,line : unsigned(8 downto 0);
	
	signal color : std_logic_vector(8 downto 0);

--Rom Teclas y Pentagrama
	signal addrTeclas: std_logic_vector (8 downto 0);
	signal bitMapTeclas: std_logic_vector (0 to 319);
	type romTypeTecla is array (0 to 239) of std_logic_vector (0 to 319);
	constant romTeclas : romTypeTecla :=(
 0=>X"00001E00000000000000000000000000000000000000000000000000000000000000000000000000", 1=>X"00001300000000000000000000000000000000000000000000000000000000000000000000000000", 2=>X"000031C0000000000000000000000000000000000000000000000000000000000000000000000000", 3=>X"00002060000000000000000000000000000000000000000000000000000000000000000000000000", 4=>X"00006020000000000000000000000000000000000000000000000000000000000000000000000000", 5=>X"0000C030000000000000000000000000000000000000000000000000000000000000000000000000", 6=>X"00018010000000000000000000000000000000000000000000000000000000000000000000000000", 7=>X"00038010000000000000000000000000000000000000000000000000000000000000000000000000", 8=>X"00070010000000000000000000000000000000000000000000000000000000000000000000000000", 9=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 10=>X"000C0030000000000000000000000000000000000000000000000000000000000000000000000000", 11=>X"001C0030000000000000000000000000000000000000000000000000000000000000000000000000", 12=>X"001C0060000000000000000000000000000000000000000000000000000000000000000000000000", 13=>X"001C00E0000000000000000000000000000000000000000000000000000000000000000000000000", 14=>X"001C00C0000000000000000000000000000000000000000000000000000000000000000000000000", 15=>X"003C0180000000000000000000000000000000000000000000000000000000000000000000000000", 16=>X"003C0380000000000000000000000000000000000000000000000000000000000000000000000000", 17=>X"003C0700000000000000000000000000000000000000000000000000000000000000000000000000", 18=>X"001C0E00000000000000000000000000000000000000000000000000000000000000000000000000", 19=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 20=>X"001C3800000000000000000000000000000000000000000000000000000000000000000000000000", 21=>X"000E7000000000000000000000000000000000000000000000000000000000000000000000000000", 22=>X"0007E000000000000000000000000000000000000000000000000000000000000000000000000000", 23=>X"0003C000000000000000000000000000000000000000000000000000000000000000000000000000", 24=>X"00038000000000000000000000000000000000000000000000000000000000000000000000000000", 25=>X"00078000000000000000000000000000000000000000000000000000000000000000000000000000", 26=>X"000EC000000000000000000000000000000000000000000000000000000000000000000000000000", 27=>X"001C6000000000000000000000000000000000000000000000000000000000000000000000000000", 28=>X"00186000000000000000000000000000000000000000000000000000000000000000000000000000", 29=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 30=>X"00387F80000000000000000000000000000000000000000000000000000000000000000000000000", 31=>X"0030F1C0000000000000000000000000000000000000000000000000000000000000000000000000", 32=>X"0061F0C0000000000000000000000000000000000000000000000000000000000000000000000000", 33=>X"00639840000000000000000000000000000000000000000000000000000000000000000000000000", 34=>X"00E71860000000000000000000000000000000000000000000000000000000000000000000000000", 35=>X"00C71860000000000000000000000000000000000000000000000000000000000000000000000000", 36=>X"00C61860C00000000000000000000000000000000000000000000000000000000000000000000000", 37=>X"00C61860C00000000000000000000000000000000000000000000000000000000000000000000000", 38=>X"00C618C0000000000000000000000000000000000000000000000000000000000000000000000000", 39=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 40=>X"00C60DC0000000000000000000000000000000000000000000000000000000000000000000000000", 41=>X"00C60D80C00000000000000000000000000000000000000000000000000000000000000000000000", 42=>X"00C60F80C00000000000000000000000000000000000000000000000000000000000000000000000", 43=>X"00C20F00000000000000000000000000000000000000000000000000000000000000000000000000", 44=>X"00C00E00000000000000000000000000000000000000000000000000000000000000000000000000", 45=>X"00603C00000000000000000000000000000000000000000000000000000000000000000000000000", 46=>X"003FF800000000000000000000000000000000000000000000000000000000000000000000000000", 47=>X"001FEC00000000000000000000000000000000000000000000000000000000000000000000000000", 48=>X"00000C00000000000000000000000000000000000000000000000000000000000000000000000000", 49=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 50=>X"00000C00000000000000000000000000000000000000000000000000000000000000000000000000", 51=>X"00001800000000000000000000000000000000000000000000000000000000000000000000000000", 52=>X"00001800000000000000000000000000000000000000000000000000000000000000000000000000", 53=>X"00001800000000000000000000000000000000000000000000000000000000000000000000000000", 54=>X"00301800000000000000000000000000000000000000000000000000000000000000000000000000", 55=>X"00FC1800000000000000000000000000000000000000000000000000000000000000000000000000", 56=>X"01FC3000000000000000000000000000000000000000000000000000000000000000000000000000", 57=>X"03883000000000000000000000000000000000000000000000000000000000000000000000000000", 58=>X"03883000000000000000000000000000000000000000000000000000000000000000000000000000", 59=>X"03003000000000000000000000000000000000000000000000000000000000000000000000000000",
 60=>X"03007000000000000000000000000000000000000000000000000000000000000000000000000000", 61=>X"0380E000000000000000000000000000000000000000000000000000000000000000000000000000", 62=>X"01FFC000000000000000000000000000000000000000000000000000000000000000000000000000", 63=>X"00FF8000000000000000000000000000000000000000000000000000000000000000000000000000", 64=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 65=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 66=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 67=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 68=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 69=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 70=>X"000FFFC0000000000000000000000000000000000000000000000000000000000000000000000000", 71=>X"001FFFF0000000000000000000000000000000000000000000000000000000000000000000000000", 72=>X"003FFFFC000000000000000000000000000000000000000000000000000000000000000000000000", 73=>X"007C01FE000000000000000000000000000000000000000000000000000000000000000000000000", 74=>X"00F0007E000000000000000000000000000000000000000000000000000000000000000000000000", 75=>X"00E0003F000000000000000000000000000000000000000000000000000000000000000000000000", 76=>X"01FF001F0C0000000000000000000000000000000000000000000000000000000000000000000000", 77=>X"01FFC01F0C0000000000000000000000000000000000000000000000000000000000000000000000", 78=>X"01FFE01F000000000000000000000000000000000000000000000000000000000000000000000000", 79=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 80=>X"01FFE01F000000000000000000000000000000000000000000000000000000000000000000000000", 81=>X"01FFE03F0C0000000000000000000000000000000000000000000000000000000000000000000000", 82=>X"01FFC07F0C0000000000000000000000000000000000000000000000000000000000000000000000", 83=>X"00FF807E000000000000000000000000000000000000000000000000000000000000000000000000", 84=>X"0000007E000000000000000000000000000000000000000000000000000000000000000000000000", 85=>X"000000FC000000000000000000000000000000000000000000000000000000000000000000000000", 86=>X"000000FC000000000000000000000000000000000000000000000000000000000000000000000000", 87=>X"000001FC000000000000000000000000000000000000000000000000000000000000000000000000", 88=>X"000003F8000000000000000000000000000000000000000000000000000000000000000000000000", 89=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 90=>X"000007E0000000000000000000000000000000000000000000000000000000000000000000000000", 91=>X"00000FC0000000000000000000000000000000000000000000000000000000000000000000000000", 92=>X"00001F80000000000000000000000000000000000000000000000000000000000000000000000000", 93=>X"00003F00000000000000000000000000000000000000000000000000000000000000000000000000", 94=>X"00007E00000000000000000000000000000000000000000000000000000000000000000000000000", 95=>X"0001FC00000000000000000000000000000000000000000000000000000000000000000000000000", 96=>X"0003F000000000000000000000000000000000000000000000000000000000000000000000000000", 97=>X"000FE000000000000000000000000000000000000000000000000000000000000000000000000000", 98=>X"001F8000000000000000000000000000000000000000000000000000000000000000000000000000", 99=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 100=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 101=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 102=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 103=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 104=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 105=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 106=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 107=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 108=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 109=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 110=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 111=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 112=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 113=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 114=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 115=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 116=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 117=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 118=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 119=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000",
 120=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 121=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 122=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 123=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 124=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 125=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 126=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 127=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 128=>X"00000000000000000000000000000000000000000000000000000000000000000000000000000000", 129=>X"FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF",
 130=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",131=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",132=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",133=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",134=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",135=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",136=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",137=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",138=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",139=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",
 140=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",141=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",142=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",143=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",144=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",145=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",146=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",147=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",148=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",149=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",
 150=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",151=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",152=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",153=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",154=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",155=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",156=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",157=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",158=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",159=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",
 160=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",161=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",162=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",163=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",164=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",165=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",166=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",167=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",168=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",169=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",
 170=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",171=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",172=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",173=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",174=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",175=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",176=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",177=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",178=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",179=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",
 180=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",181=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",182=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",183=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",184=>X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FFF00FFFF7FFFF8",185=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",186=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",187=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",188=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",189=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",
 190=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",191=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",192=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",193=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",194=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",195=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",196=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",197=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",198=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",199=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",
 200=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",201=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",202=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",203=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",204=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",205=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",206=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",207=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",208=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",209=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",
 210=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",211=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",212=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",213=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",214=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",215=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",216=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",217=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",218=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",219=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",
 220=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",221=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",222=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",223=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",224=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",225=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",226=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",227=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",228=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",229=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",
 230=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",231=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",232=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",233=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",234=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",235=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",236=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",237=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",238=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8",239=>X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8"
 );


--0001 1111 1111 1111 1111 1110 000 0 0000 1111 1111 0000 0 000 0111 1111 1111 1111 1 0 11 1111 1111 1111 1100 00 0 0 0001 1111 1111 1110 000 0 0000 1111 1111 1111 0000 0 000 0111 1111 1111 1111 0 1 11 1111 1111 1111 1100 00 0 0 0001 1111 1111 1110 000 0 0000 1111 1111 1111 1111 0 111 1111 1111 1111 1000 0 0 00 0011 1111 1111 1100 00 0 0 0001 1111 1111 1111 000 0 0000 1111 1111 1111 1111 0 111 1111 1111 1111 1111 1000
--1    F     F    F    F    E    0      0    F    F    0     0    7    F    F   F      B    F     F    F   C      0     1    F    F    E     0    0    F    F    F    0     0    7    F    F    F     7     F    F    F    C      0    1    F    F    E     0    0    F    F    F    F    7     F    F    F    8      0     3   F    F    C      0    1   F     F    F     0    0    F    F    F    F    7     F    F    F    F    8
 --  
--
--1     F     F    F   F    F    E      F   F    F    F     7     F    F   F     F    B      F    F    F    F    B     F     F    F    F    E     F    F    F   F     F     7   F    F     F    F    7      F    F    F    F    B     F     F    F    F    E     F    F    F    F    F     7   F     F    F    F    7      F    F    F    F    B      F    F    F    F   E      F   F     F    F    F     7   F     F    F    F   8 
--0001 1111 1111 1111 1111 1111 111 0 1111 1111 1111 1111 0 111 1111 1111 1111 1111 1 0 11 1111 1111 1111 1111 11 0 1 1111 1111 1111 1111 111 0 1111 1111 1111 1111 1111 0 111 1111 1111 1111 1111 0 1 11 1111 1111 1111 1111 11 0 1 1111 1111 1111 1111 111 0 1111 1111 1111 1111 1111 0 111 1111 1111 1111 1111 0 1 11 1111 1111 1111 1111 11 0 1 1111 1111 1111 1111 111 0 1111 1111 1111 1111 1111 0 111 1111 1111 1111 1111 1000
--			DOF										REF								MIF								FF										SolF								LAF										SIF					DO											RE										Mi						FA											Sol								LA										Si							Do
--
--X"1FFFFE00FF007FF803FFC01FFE00FFF007FF803FFC01FFE00FFF007FF803FFC01FFE00FFF007FFF8"
--Parte Superior
--X"1FFFFE00FF007FFFBFFFC01FFE00FFF007FFF7FFFC01FFE00FFFF7FFF803FFC01FF700FFFF7FFFF8"
--Parte Inferior
--X"1FFFFFEFFFF7FFFFBFFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF7FFFFBFFFFEFFFFF7FFFF8"

--Rom Nota
signal addrNota: std_logic_vector (4 downto 0);
	signal bitMapNota: std_logic_vector (0 to 15);
	type romTypeNota is array (0 to 8) of std_logic_vector (0 to 15);
	signal romNota : romTypeNota :=(0=>X"0000", 1=>X"0000",2=>X"0180", 3=>X"03C0", 4=>X"07E0", 5=>X"07E0", 6=>X"03C0", 7=>X"0180", 8=>X"0000");

--Rom Nota Alterada
signal addrNotaAlt: std_logic_vector (4 downto 0);
	signal bitMapNotaAlt: std_logic_vector (0 to 15);
	signal romNotaAlt : romTypeNota :=(0=>X"0008", 1=>X"000F",2=>X"0189", 3=>X"03CF", 4=>X"07E0", 5=>X"07E0", 6=>X"03C0", 7=>X"0180", 8=>X"0000");


begin

	
  screenInteface: vgaInterface
  generic map ( FREQ => 50_000, SYNCDELAY => 0 )
  port map ( rst_n => rst_n, clk => clk, line => lineAux, pixel => pixelAux, R => color(8 downto 6), G => color(5 downto 3), B => color(2 downto 0), hSync => hSync, vSync => vSync, RGB => RGB );
----------------------------------------------------------------------------------------------------------------------------------------------------------------


	selectColor:
	process(Pentagramas,Notas,line,colorVerde,colorAzul)
	begin
		if Pentagramas='1' or Notas='1' then
		  if line=129 then
			color<="101000000";
		  elsif colorVerde='1' then
            color<="000101000";
        else
            color<=(others=>'1');
		  end if;
		else
		  if colorAzul='1' then
            color<="000000100";
		  else
			color<=(others=>'0');
		  end if;
		end if;
	end process;

	pixel <= unsigned(pixelAux(9 downto 1));
	line <= unsigned(lineAux(9 downto 1));
	
	Pentagramas <= bitMapTeclas(to_integer(pixel));
						
	addrTeclas<=std_logic_vector(line);	
	
	romTeclitas : process(clk)
	begin
      if rising_edge(clk) then
			bitMapTeclas <=romTeclas(to_integer(unsigned(addrTeclas)));
		end if;
	end process;


	colorAzul<= '1' when (teclaPulsadaPintar(1)='1' or teclaPulsadaPintar(3)='1' or teclaPulsadaPintar(6)='1'or teclaPulsadaPintar(8)='1' or teclaPulsadaPintar(10)='1' or 
								teclaPulsadaPintar(13)='1' or teclaPulsadaPintar(15)='1' or teclaPulsadaPintar(18)='1' or teclaPulsadaPintar(20)='1' or teclaPulsadaPintar(22)='1'
								) else '0';
	--rebF
	teclaPulsadaPintar(1)<= '1' when (pixel>=23 and pixel<=31 and line>129 and line<185 and teclaPulsada(1)='1') else '0';
	--mibF
	teclaPulsadaPintar(3)<= '1' when (pixel>=40 and pixel<=48 and line>129 and line<185 and teclaPulsada(3)='1') else '0';
	--solbF
	teclaPulsadaPintar(6)<= '1' when (pixel>=82 and pixel<=90 and line>129 and line<185 and teclaPulsada(6)='1') else '0';
	--labF
	teclaPulsadaPintar(8)<= '1' when (pixel>=103 and pixel<=111 and line>129 and line<185 and teclaPulsada(8)='1') else '0';	
	--sibF
	teclaPulsadaPintar(10)<= '1' when (pixel>=124 and pixel<=132 and line>129 and line<185 and teclaPulsada(10)='1') else '0';
	--reb
	teclaPulsadaPintar(13)<= '1' when (pixel>=166 and pixel<=174 and line>129 and line<185 and teclaPulsada(13)='1') else '0';
	--mib
	teclaPulsadaPintar(15)<= '1' when (pixel>=187 and pixel<=195 and line>129 and line<185 and teclaPulsada(15)='1') else '0';
	--solb
	teclaPulsadaPintar(18)<= '1' when (pixel>=229 and pixel<=237 and line>129 and line<185 and teclaPulsada(18)='1') else '0';
	--lab
	teclaPulsadaPintar(20)<= '1' when (pixel>=250 and pixel<=258 and line>129 and line<185 and teclaPulsada(20)='1') else '0';
	--sib
	teclaPulsadaPintar(22)<= '1' when (pixel>=272 and pixel<=279 and line>129 and line<185 and teclaPulsada(22)='1') else '0';
	
	
	
	colorVerde<= '1' when (teclaPulsadaPintar(0)='1' or teclaPulsadaPintar(2)='1' or teclaPulsadaPintar(4)='1'or teclaPulsadaPintar(5)='1' or teclaPulsadaPintar(7)='1' or teclaPulsadaPintar(9)='1' or teclaPulsadaPintar(11)='1' or 
								  teclaPulsadaPintar(12)='1' or teclaPulsadaPintar(14)='1' or teclaPulsadaPintar(16)='1' or teclaPulsadaPintar(17)='1' or teclaPulsadaPintar(19)='1' or teclaPulsadaPintar(21)='1' or teclaPulsadaPintar(23)='1' or teclaPulsadaPintar(24)='1'
								  ) else '0';
	
	--DoF
	teclaPulsadaPintar(0)<= '1' when ( (pixel>=3 and pixel<=22 and line>129 and line<185) or (pixel>=3 and pixel<=26 and line>=185 and line<240) )and teclaPulsada(0)='1'  else '0';
	--ReF
	teclaPulsadaPintar(2)<= '1' when ( (pixel>=32 and pixel<=39 and line>129 and line<185) or (pixel>=28 and pixel<=43 and line>=185 and line<240) )and teclaPulsada(2)='1'  else '0';
	--MiF
	teclaPulsadaPintar(4)<= '1' when ( (pixel>=49 and pixel<=64 and line>129 and line<240) or (pixel>=45 and pixel<=64 and line>=185 and line<240) )and teclaPulsada(4)='1'  else '0';
	--FaF
	teclaPulsadaPintar(5)<= '1' when ((pixel>=66 and pixel<=81 and line>129 and line<185) or (pixel>=66 and pixel<=85 and line>=185 and line<240) ) and teclaPulsada(5)='1'  else '0';
	--SolF
	teclaPulsadaPintar(7)<= '1' when ( (pixel>=91 and pixel<=102 and line>129 and line<185) or (pixel>=86 and pixel<=106 and line>=185 and line<240) )and teclaPulsada(7)='1'  else '0';
	--LaF
	teclaPulsadaPintar(9)<= '1' when ( (pixel>=112 and pixel<=124 and line>129 and line<185) or (pixel>=108 and pixel<=127 and line>=185 and line<240) )and teclaPulsada(9)='1'  else '0';
	--SiF
	teclaPulsadaPintar(11)<= '1' when ((pixel>=133 and pixel<=147 and line>129 and line<240) or (pixel>=129 and pixel<=147 and line>=185 and line<240) )  and teclaPulsada(11)='1'  else '0';
	--Do
	teclaPulsadaPintar(12)<= '1' when ( (pixel>=149 and pixel<=165 and line>129 and line<185) or (pixel>=149 and pixel<=169 and line>=185 and line<240) )and teclaPulsada(12)='1'  else '0';
	--Re
	teclaPulsadaPintar(14)<= '1' when ( (pixel>=175 and pixel<=186 and line>129 and line<185) or (pixel>=170 and pixel<=190 and line>=185 and line<240) )and teclaPulsada(14)='1'  else '0';
	--Mi
	teclaPulsadaPintar(16)<= '1' when ( (pixel>=196 and pixel<=211 and line>129 and line<185) or (pixel>=192 and pixel<=211 and line>=185 and line<240) )and teclaPulsada(16)='1'  else '0';
	--Fa
	teclaPulsadaPintar(17)<= '1' when ( (pixel>=213 and pixel<=228 and line>129 and line<185) or (pixel>=213 and pixel<=232 and line>=185 and line<240) )and teclaPulsada(17)='1'  else '0';
	--Sol
	teclaPulsadaPintar(19)<= '1' when ( (pixel>=237 and pixel<=249 and line>129 and line<185) or (pixel>=233 and pixel<=253 and line>=185 and line<240) )and teclaPulsada(19)='1'  else '0';
	--La
	teclaPulsadaPintar(21)<= '1' when ( (pixel>=259 and pixel<=271 and line>129 and line<185) or (pixel>=254 and pixel<=274 and line>=185 and line<240) )and teclaPulsada(21)='1'  else '0';
	--Si
	teclaPulsadaPintar(23)<= '1' when ( (pixel>=280 and pixel<=295 and line>129 and line<185) or (pixel>=276 and pixel<=295 and line>=185 and line<240) )and teclaPulsada(23)='1'  else '0';
	--Do1
	teclaPulsadaPintar(24)<= '1' when (pixel>=297 and pixel<=316 and line>129 and line<240)and teclaPulsada(24)='1'  else '0';

--Pintar Notas

	nota(0)<= '1' when line>89 and line<99 and pixel>=25 and pixel<=40  else '0'; --Do FA
	nota(1)<= '1' when line>83 and line<93 and pixel>=38 and pixel<=53  else '0'; --reb y re FA
	nota(2)<= '1' when line>79 and line<89 and pixel>=54 and pixel<=69 else '0'; --mi y mib FA
	nota(3)<= '1' when line>73 and line<83 and pixel>=70 and pixel<=85 else '0'; --Fa FA
	nota(4)<= '1' when line>69 and line<79 and pixel>=86 and pixel<=101 else '0'; --Sol FA y Solb FA
	nota(5)<= '1' when line>63 and line<73 and pixel>=102 and pixel<=117 else '0'; --La y Lab FA
	nota(6)<= '1' when line>59 and line<69 and pixel>=118 and pixel<=133	else '0'; --Si y Sib FA
	nota(7)<= '1' when line>53 and line<63 and pixel>=134 and pixel<=149 else '0'; --Do
	nota(8)<= '1' when line>49 and line<59 and pixel>=150 and pixel<=165 else '0'; --Re y reB
	nota(9)<= '1' when line>43 and line<53 and pixel>=166 and pixel<=181 else '0'; --Mi y mib
	nota(10)<= '1' when line>39 and line<49 and pixel>=182 and pixel<=196 else '0'; --Fa
	nota(11)<= '1' when line>33 and line<43 and pixel>=197 and pixel<=212 else '0'; --Sol y solb
	nota(12)<= '1' when line>29 and line<39 and pixel>=213 and pixel<=228 else '0'; --La y lab
	nota(13)<= '1' when line>23 and line<33 and pixel>=229 and pixel<=244 else '0'; --Si y sib
	nota(14)<= '1' when line>19 and line<29 and pixel>=245 and pixel<=260 else '0'; --Do1



	selectAddrNota : process(line,nota)
	begin
		addrNota<="01000";
		addrNotaAlt<="01000";
		dir <= (others => '0');
	   if nota(0)='1' then
			dir<=std_logic_vector(line-90); --Do F
			addrNota<=dir(4 downto 0);
	   elsif nota(1)='1' then
			dir<=std_logic_vector(line-84);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Re F
	   elsif nota(2)='1' then
			dir<=std_logic_vector(line-80);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Mi F
	   elsif nota(3)='1' then
			dir<=std_logic_vector(line-74); --Fa F
			addrNota<=dir(4 downto 0);
	  elsif nota(4)='1' then 
			dir<=std_logic_vector(line-70);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Sol F
	  elsif nota(5)='1' then
			dir<=std_logic_vector(line-64);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --La F			
	  elsif nota(6)='1' then
			dir<=std_logic_vector(line-60); 
			addrNota<=dir(4 downto 0);--Si F
			addrNotaAlt<=dir(4 downto 0);--Sib F
	  elsif nota(7)='1' then
			dir<=std_logic_vector(line-54); --Do 
			addrNota<=dir(4 downto 0);
	  elsif nota(8)='1' then
			dir<=std_logic_vector(line-50);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Re      
	  elsif nota(9)='1' then
			dir<=std_logic_vector(line-44);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Mi   
	  elsif nota(10)='1' then
			dir<=std_logic_vector(line-40); --Fa   
			addrNota<=dir(4 downto 0);
	  elsif nota(11)='1' then
			dir<=std_logic_vector(line-34);  
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Sol   
	  elsif nota(12)='1' then
			dir<=std_logic_vector(line-30);
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --La   
	  elsif nota(13)='1' then
  			dir<=std_logic_vector(line-24); 
			addrNotaAlt<=dir(4 downto 0);
			addrNota<=dir(4 downto 0); --Si   
	  elsif nota(14)='1' then
			dir<=std_logic_vector(line-20); --Do1   
			addrNota<=dir(4 downto 0);
		end if;
	end process;



romNotita : process(clk)
	begin
      if rising_edge(clk) then
			bitMapNota <=romNota(to_integer(unsigned(addrNota)));
		end if;
	end process;

romNotaAlterada : process(clk)
	begin
      if rising_edge(clk) then
			bitMapNotaALt <=romNotaAlt(to_integer(unsigned(addrNotaAlt)));
		end if;
	end process;



	Notas<= '1' when (  notaPintar(0)='1'  or  notaPintar(1)='1' or notaPintar(2)='1' or notaPintar(3)='1' or notaPintar(4)='1' or notaPintar(5)='1' or notaPintar(6)='1' or notaPintar(7)='1' or notaPintar(8)='1' or notaPintar(9)='1' or notaPintar(10)='1' or notaPintar(11)='1' or notaPintar(12)='1' or notaPintar(13)='1' 
					or notaPintar(14)='1' or notaPintar(15)='1' or notaPintar(16)='1' or notaPintar(17)='1' or notaPintar(18)='1' or notaPintar(19)='1' or notaPintar(20)='1' or notaPintar(21)='1' or notaPintar(22)='1' or notaPintar(23)='1' or notaPintar(24)='1' 
					)else'0';

	--DoF
	notaPintar(0)<= '1' when  (nota(0)='1' and bitMapNota(to_integer(pixel-25))='1') and teclaPulsada(0)='1'  else '0';
	--ReF
	notaPintar(2)<= '1' when  (nota(1)='1' and bitMapNota(to_integer(pixel-38))='1' ) and teclaPulsada(2)='1'  else '0';
	--MiF
	notaPintar(4)<= '1' when (nota(2)='1' and bitMapNota(to_integer(pixel-54))='1'  )and teclaPulsada(4)='1'  else '0';
	--FaF
	notaPintar(5)<= '1' when (nota(3)='1' and bitMapNota(to_integer(pixel-70))='1' ) and teclaPulsada(5)='1'  else '0';
	--SolF
	notaPintar(7)<= '1' when ( nota(4)='1' and bitMapNota(to_integer(pixel-86))='1' )and teclaPulsada(7)='1'  else '0';
	--LaF
	notaPintar(9)<= '1' when ( nota(5)='1' and bitMapNota(to_integer(pixel-102))='1')and teclaPulsada(9)='1'  else '0';
	--SiF
	notaPintar(11)<= '1' when (nota(6)='1' and bitMapNota(to_integer(pixel-118))='1' )  and teclaPulsada(11)='1'  else '0';
	--Do
	notaPintar(12)<= '1' when ( nota(7)='1' and ( ( pixel>=135 and pixel<=148 and (line=59 or line=58) ) or bitMapNota(to_integer(pixel-134))='1') )and teclaPulsada(12)='1'  else '0';
	--Re
	notaPintar(14)<= '1' when ( nota(8)='1' and ( bitMapNota(to_integer(pixel-150))='1'))and teclaPulsada(14)='1'  else '0';
	--Mi
	notaPintar(16)<= '1' when ( nota(9)='1' and ( bitMapNota(to_integer(pixel-166))='1'))and teclaPulsada(16)='1'  else '0';
	--Fa
	notaPintar(17)<= '1' when ( nota(10)='1' and ( bitMapNota(to_integer(pixel-182))='1') )and teclaPulsada(17)='1'  else '0';
	--Sol
	notaPintar(19)<= '1' when ( nota(11)='1' and ( bitMapNota(to_integer(pixel-197))='1'))and teclaPulsada(19)='1'  else '0';
	--La
	notaPintar(21)<= '1' when ( nota(12)='1' and ( bitMapNota(to_integer(pixel-213))='1'))and teclaPulsada(21)='1'  else '0';
	--Si
	notaPintar(23)<= '1' when ( nota(13)='1' and ( bitMapNota(to_integer(pixel-229))='1'))and teclaPulsada(23)='1'  else '0';
	--Do1
	notaPintar(24)<= '1' when (nota(14)='1' and ( bitMapNota(to_integer(pixel-245))='1'))and teclaPulsada(24)='1'  else '0';

	--rebF
	notaPintar(1)<= '1' when (nota(1)='1' and  bitMapNotaAlt(to_integer(pixel-38))='1' and teclaPulsada(1)='1') else '0';
	--mibF
	notaPintar(3)<= '1' when ( nota(2)='1' and bitMapNotaAlt(to_integer(pixel-54))='1' and teclaPulsada(3)='1') else '0';
	--solbF
	notaPintar(6)<= '1' when (nota(4)='1' and bitMapNotaAlt(to_integer(pixel-86))='1' and teclaPulsada(6)='1') else '0';
	--labF
	notaPintar(8)<= '1' when ( nota(5)='1' and  bitMapNotaAlt(to_integer(pixel-102))='1' and teclaPulsada(8)='1') else '0';	
	--sibF
	notaPintar(10)<= '1' when ( nota(6)='1' and  bitMapNotaAlt(to_integer(pixel-118))='1' and teclaPulsada(10)='1') else '0';
	--reb
	notaPintar(13)<= '1' when (nota(8)='1' and  bitMapNotaAlt(to_integer(pixel-150))='1' and teclaPulsada(13)='1') else '0';
	--mib
	notaPintar(15)<= '1' when (nota(9)='1' and  bitMapNotaAlt(to_integer(pixel-166))='1' and teclaPulsada(15)='1') else '0';
	--solb
	notaPintar(18)<= '1' when (nota(11)='1' and  bitMapNotaAlt(to_integer(pixel-197))='1' and teclaPulsada(18)='1') else '0';
	--lab
	notaPintar(20)<= '1' when (nota(12)='1' and  bitMapNotaAlt(to_integer(pixel-213))='1' and teclaPulsada(20)='1') else '0';
	--sib
	notaPintar(22)<= '1' when (nota(13)='1' and  bitMapNotaAlt(to_integer(pixel-229))='1' and teclaPulsada(22)='1') else '0';	 

end Behavioral;

